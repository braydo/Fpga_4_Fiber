`timescale 1ns/100ps

module MPD (
	inout [31:0] VME_DATA,
	inout [31:0] VME_ADDR,
	input [5:0] VME_AM,
	input [5:0] VME_GA,
	input VME_WRITEb,
	input VME_DS0b,
	input VME_DS1b,
	input VME_ASb,
	input VME_IACKb,
	input VME_IACKINb,
	output VME_IACKOUTb,
	output VME_DTACKb,
	output VME_BERRb,
	output VME_RETRYb,

	output APV_CLOCK, output APV_TRIGGER, output APV_RESET,
	output I2C_SCL, inout I2C_SDA,

	input [1:0] USER_IN, output [1:0] USER_OUT,	// USER_IN[0] = trigger, USER_IN[1] = sync
	input CLK_FRONT,

	output GXB_TX, input GXB_RX, input GXB_PRESENT, input GXB_RX_LOS,

//	input [1:0] ADC_PATTERN,	// Debug: simulate APV frames 0 = ADC_Deskew, 1 = ADC_Sync, 2 = APV_SYNC, 3 = APV_FRAME
	input APV_SAMPLE_MODE,	// 0 = 3 samples, 1 = 1 sample
	output FIBER_LINK_READY
);

parameter master_ck_period = 25;
parameter master_ck_half_period = master_ck_period / 2;
parameter master_ck_hold  = 1;	// data hold time

parameter fast_ck_period = 16;
parameter fast_ck_half_period = fast_ck_period / 2;

parameter gxb_ck_period = 16;
parameter gxb_ck_half_period = gxb_ck_period / 2;

reg Master_clock, Master_resetB;
wire adc_lclk1, adc_lclk2, adc_ck1, adc_ck2, adc_conv_ck;
wire [15:0] adc_data;
wire [31:0] vme_data_x, vme_addr_x;
wire vme_dtackB_x, vme_berrB_x, vme_retryB_x;
wire Sdram_ck, Sdram_ckB, Sdram_rasB, Sdram_casB, Sdram_weB, Sdram_dm, Sdram_odt;
wire Sdram_csB, Sdram_cke;
wire [2:0] Sdram_ba;
wire [13:0] Sdram_addr;
tri1 [7:0] Sdram_dq;
tri1 [7:1] vme_irqB;
tri1 Sdram_dqsN;	// same as wire
tri0 Sdram_dqs;		// same as wire
reg trig_pulse;
reg fast_clock, gxb_clock;
wire [3:0] leds;


assign FIBER_LINK_READY = leds[3];

BidirBuf #(32) Abuf(.A(vme_addr_x), .B(VME_ADDR), .OEb(vme_aoeB), .DIR(vme_adir));
BidirBuf #(32) Dbuf(.A(vme_data_x), .B(VME_DATA), .OEb(vme_doeB), .DIR(vme_ddir));
BidirBuf #(1) Dtack_buf(.A(vme_dtackB_x), .B(VME_DTACKb), .OEb(~vme_dtack_en), .DIR(1'b1));
BidirBuf #(1) Berr_buf(.A(vme_berrB_x), .B(VME_BERRb), .OEb(~vme_berr_en), .DIR(1'b1));
BidirBuf #(1) Retry_buf(.A(vme_retryB_x), .B(VME_RETRYb), .OEb(~vme_retry_en), .DIR(1'b1));

Fpga Dut(
	.MASTER_RESETb(Master_resetB), .MASTER_CLOCK(Master_clock), .MASTER_CLOCK2(CLK_FRONT),

	.VME_D(vme_data_x), .VME_A(vme_addr_x), .VME_AM(VME_AM), .VME_GA(VME_GA),
	.VME_WRITEb(VME_WRITEb), .VME_DS0b(VME_DS0b), .VME_DS1b(VME_DS1b), .VME_ASb(VME_ASb),
	.VME_IACKb(VME_IACKb), .VME_IACKINb(VME_IACKINb), .VME_IACKOUTb(VME_IACKOUTb),
	.VME_DTACKb(vme_dtackB_x), .VME_BERRb(vme_berrB_x), .VME_RETRYb(vme_retryB_x),
	.VME_IRQ(vme_irqB), .VME_ADIR(vme_adir), .VME_AOEb(vme_aoeB),
	.VME_DDIR(vme_ddir), .VME_DOEb(vme_doeB),
	.VME_DTACK_EN(vme_dtack_en), .VME_BERR_EN(vme_berr_en), .VME_RETRY_EN(vme_retry_en),
	.VME_LIIb(), .VME_LIOb(),

	.ADC_DATA(adc_data), .ADC_RESETb(adc_resetB),
	.ADC_CS1b(adc_cs1B), .ADC_CS2b(adc_cs2B), .ADC_SCLK(adc_sclk), .ADC_SDA(adc_sda),
	.ADC_LCLK1(adc_lclk1), .ADC_LCLK2(adc_lclk2), .ADC_FRAME_CK1(adc_ck1), .ADC_FRAME_CK2(adc_ck2),
	.ADC_CONV_CK1(adc_conv_ck),

	.APV_CLOCK(APV_CLOCK), .APV_TRIGGER(APV_TRIGGER), .APV_RESET(APV_RESET),

	.I2C_SCL(I2C_SCL), .I2C_SDA_IN(I2C_SDA), .I2C_SDA_OUT(I2C_SDA),

	.USER_IN_TTL(USER_IN), .USER_IN_NIM(~USER_IN), .USER_OUT(USER_OUT), .SEL_OUT(),

	.MII_25MHZ_CLOCK(), .MII_MDC(), .MII_MDIO(),
	.MII_TX_CLK(), .MII_TX_EN(), .MII_TXD(),
	.MII_RX_CLK(), .MII_RX_DV(), .MII_RX_ER(), .MII_RXD(),
	.MII_CRS(), .MII_COL(), .MII_RESETb(),

	.SDRAM_A(Sdram_addr), .SDRAM_BA(Sdram_ba), .SDRAM_CASb(Sdram_casB), .SDRAM_CKE(Sdram_cke),
	.SDRAM_CSb(Sdram_csB), .SDRAM_DM(Sdram_dm), .SDRAM_RASb(Sdram_rasB), .SDRAM_WEb(Sdram_weB),
	.SDRAM_CK(Sdram_ck), .SDRAM_CKb(Sdram_ckB), .SDRAM_DQ(Sdram_dq), .SDRAM_DQS(Sdram_dqs), .SDRAM_ODT(Sdram_odt),

	.SD_DAT2(), .SD_DAT1(), .SD_DAT0(), .SD_DETECT(), .SD_CD(), .SD_CMD(), .SD_CLK(),
	
	.READ1(), .READ_CLK1(),	.READ2(), .READ_CLK2(),

	.LED(leds), .SWITCH(4'b1111),

	.GXB_TX(GXB_TX), .GXB_RX(GXB_RX), .GXB_PRESENT(GXB_PRESENT),
	.GXB_TX_DISABLE(), .GXB_RX_LOS(GXB_RX_LOS), .GXB_CK(gxb_clock),

	.TOKEN_OUT_P0(), .TOKEN_OUT_P2(), .TOKEN_IN_P0(1'b0), .TOKEN_IN_P2(1'b0),
	.TRIG_OUT(), .BUSY_OUT(), .SD_LINK_OUT(),
	.TRIG1_IN(1'b0), .TRIG2_IN(1'b0), .SYNC_IN(1'b0), .STATBIT_A_IN(1'b0), .STATBIT_B_IN(1'b0), .CLK_IN_P0(fast_clock),
	.STATBIT_A_OUT(),

	.SPARE1(), .SPARE2(), .SPARE3(),
	
	.SPARE33(),
	.SPARE25(),
	.SPARE_CLK_LVDS(), .SPARE_CLK_TTL()

);
/*
// This is MICRON model
ddr2 Sdram0(.ck(Sdram_ck), .ck_n(Sdram_ckB), .cke(Sdram_cke), .cs_n(Sdram_csB),
	.ras_n(Sdram_rasB), .cas_n(Sdram_casB), .we_n(Sdram_weB), .ba(Sdram_ba), .addr(Sdram_addr),
	.dm_rdqs(Sdram_dm), .dq(Sdram_dq), .dqs(Sdram_dqs), .odt(Sdram_odt), .dqs_n(Sdram_dqsN), .rdqs_n());
*/

// This model is generated by DDR Controller MegaWizard
Ddr2SdramIf_full_mem_model Sdram0(
                                    // inputs:
                                     .mem_addr(Sdram_addr),
                                     .mem_ba(Sdram_ba),
                                     .mem_cas_n(Sdram_casB),
                                     .mem_cke(Sdram_cke),
                                     .mem_clk(Sdram_ck),
                                     .mem_clk_n(Sdram_ckB),
                                     .mem_cs_n(Sdram_csB),
                                     .mem_dm(Sdram_dm),
                                     .mem_odt(Sdram_odt),
                                     .mem_ras_n(Sdram_rasB),
                                     .mem_we_n(Sdram_weB),

                                    // outputs:
                                     .global_reset_n(),
                                     .mem_dq(Sdram_dq),
                                     .mem_dqs(Sdram_dqs),
                                     .mem_dqs_n(Sdram_dqsN)
                                  );
	
ads5281_apv ADC1(.APV_TRIGGER(APV_TRIGGER), .APV_MODE(APV_SAMPLE_MODE), .CLK(adc_conv_ck),
	.LCLK(adc_lclk1), .ADCLK(adc_ck1), .OUT18(adc_data[7:0]));
ads5281_apv ADC2(.APV_TRIGGER(APV_TRIGGER), .APV_MODE(APV_SAMPLE_MODE), .CLK(adc_conv_ck),
	.LCLK(adc_lclk2), .ADCLK(adc_ck2), .OUT18(adc_data[15:8]));
defparam ADC1.data_file_prefix = "/home/braydo/Projects/fe_fw/Simulation/aldec/default/testbench/mpd_data/apv_data0_";
defparam ADC2.data_file_prefix = "/home/braydo/Projects/fe_fw/Simulation/aldec/default/testbench/mpd_data/apv_data1_";

  // Clock generator: free running
  initial
  begin
    #(master_ck_period-master_ck_hold)	Master_clock <= ~Master_clock;
    forever
      #master_ck_half_period	Master_clock <= ~Master_clock;
  end

  always
	  #fast_ck_half_period fast_clock = ~fast_clock;

  always
	  #gxb_ck_half_period gxb_clock = ~gxb_clock;

  initial	// Power UP Reset
  begin
	     Master_resetB = 1;
	     Master_clock = 0;
	     fast_clock = 0;
	     gxb_clock = 0;
	#1000 Master_resetB = 0;
	#100 Master_resetB = 1;
  end

endmodule

